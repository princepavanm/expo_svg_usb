`include "usbf_crc16.v"
`include "usbf_crc5.v"
`include "usbf_defines.v"

`include "usbf_utmi_ls.v"
`include "usbf_utmi_if.v"

`include "usbf_idma.v"
`include "usbf_pa.v"
`include "usbf_pd.v"
`include "usbf_pe.v"
`include "usbf_pl.v"

`include "usbf_mem_arb.v"

`include "usbf_ep_rf.v"
//`include "usbf_ep_rf_dummy.v"
`include "usbf_rf.v"

`include "usbf_wb.v"

`include "usbf_top.v"
