//List of Include Files

  `include "usb_base_test.sv"

