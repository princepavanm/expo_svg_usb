///////////////////////////////////////////////////////////////////////////////////////////////////
//      Company:  Expolog Technologies.                                                          //
//           Copyright (c) 2023 by Expolog Technologies, Inc. All rights reserved.               //
//                                                                                               //
//      Engineer          :  ANGAPPAN, MOHAMMED_KHADEER, LOKESH, MADHURA.                        //
//      Revision Tag      :  06/10/2023                                                          //                                                   
//      Project Name      :  USB 3.1                                                             //
//      Component Name    :  Sequence_list                                                       //
//      Description       :  All sequence files are listed.                                      // 
//                                                                                               //
//                                                                                               //
//                                                                                               // 
//      Additional Comments:                                                                     //
//                                                                                               //
///////////////////////////////////////////////////////////////////////////////////////////////////

  //List of Include Files

  `include "reset_sequence.sv"
  `include "mid_reset_seq.sv"
  `include "debug_sof_seq.sv"
  `include "usb_base_seq.sv"
  `include "speed_neg_hs_seq.sv"
  `include "phy_rx_seq.sv"
  `include "token_in_seq.sv"
`include "token_out_ep1_seq.sv"
