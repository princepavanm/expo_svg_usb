//List of Include Files

  `include "utmi_base_seq.sv"




