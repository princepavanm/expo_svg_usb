//List of Include Files

  `include "utmi_base_seq.sv"

  `include "utmi_speed_neg_seq.sv"
  `include "utmi_fs_speed_neg_seq.sv"


