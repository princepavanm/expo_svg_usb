//List of Include Files

  `include "usb_base_seq.sv"
  `include "reset_sequence.sv"

