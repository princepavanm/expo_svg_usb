/* PROJECT NAME: USB 
*/
