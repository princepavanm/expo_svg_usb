///////////////////////////////////////////////////////////////////////////////////////////////////
//      Company:  Expolog Technologies.                                                          //
//           Copyright (c) 2023 by Expolog Technologies, Inc. All rights reserved.               //
//                                                                                               //
//      Engineer          :  ANGAPPAN, MOHAMMED_KHADEER, LOKESH, MADHURA.                        //
//      Revision tag      :  06/10/2023                                                          //                                                   
//      Project Name      :  USB 3.1                                                             //
//      component name    :  Sequence_list                                                       //
//      Description       :  all sequence files are listed.                                      //   
//     Additional Comments:                                                                      //
//                                                                                               //
///////////////////////////////////////////////////////////////////////////////////////////////////

//List of Include Files

  `include "reset_sequence.sv"
  `include "usb_base_seq.sv"
  `include "phy_rx_seq.sv"

