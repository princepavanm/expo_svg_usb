//List of Include Files

  `include "reset_intf.sv"
  `include "wb_agent_intf.sv"
  `include "utmi_agent_intf.sv"
  `include "sram_agent_intf.sv"

  `include "reset_tx.sv"
  `include "reset_driver.sv"
  //`include "reset_sqr.sv"
  `include "reset_agent.sv"

  `include "wb_agent_tx.sv"
  `include "wb_agent_drv.sv"
  `include "wb_agent_sqr.sv"
  `include "wb_agent_cov.sv"
  `include "wb_agent_mon.sv"
  `include "wb_agent.sv"

  `include "utmi_agent_tx.sv"
  `include "utmi_agent_drv.sv"
  `include "utmi_agent_sqr.sv"
  `include "utmi_agent_cov.sv"
  `include "utmi_agent_mon.sv"
  `include "utmi_agent.sv"

  `include "sram_agent_tx.sv"
  `include "sram_agent_drv.sv"
  `include "sram_agent_sqr.sv"
  `include "sram_agent_cov.sv"
  `include "sram_agent_mon.sv"
  `include "sram_agent.sv"

  `include "virtual_sqr.sv"

// Sequence List
  `include "../seqs/sequence_list.sv"
  `include "env.sv"

// Test List
  `include "../tests/test_list.sv"
