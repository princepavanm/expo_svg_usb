//List of Include Files

  `include "usb_base_test.sv"
  `include "usb_reg_reset_read_test.sv"
  `include "usb_reg_write_read_test.sv"
  `include "usb_reg_reset_read_reg_model_test.sv"
  `include "usb_reg_write_read_reg_model_test.sv"
  `include "utmi_speed_neg_test.sv"
  `include "utmi_fs_speed_neg_test.sv"

