//List of Include Files

  `include "wb_base_seq.sv"
  `include "reset_sequence.sv"
  `include "wb_reg_reset_read_seq.sv"
  `include "wb_reg_write_read_seq.sv"
  `include "wb_reg_reset_read_reg_model_seq.sv"
  `include "wb_reg_write_read_reg_model_seq.sv"
  `include "wb_usb_config_seq.sv"
  `include "wb_intr_handling_seq.sv"

