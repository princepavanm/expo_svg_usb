///////////////////////////////////////////////////////////////////////////////////////////////////
//      Company:  Expolog Technologies.                                                          //
//           Copyright (c) 2023 by Expolog Technologies, Inc. All rights reserved.               //
//                                                                                               //
//      Engineer          :  ANGAPPAN, MOHAMMED_KHADEER, LOKESH, MADHURA.                        //
//      Revision Tag      :  06/10/2023                                                          //
//      Module Name       :  Test_list                                                           //
//      Project Name      :  USB 3.1                                                             //
//      Component Name    :  test_list                                                           //
//      Description       :  In this file all test bench files are included.                     //
//                                                                                               //
//                                                                                               //
//     Additional Comments:                                                                      //
//                                                                                               //
///////////////////////////////////////////////////////////////////////////////////////////////////

  //List of Include Files
  	`include "usb_base_test.sv"
	`include "usb_mid_reset_test.sv"
   	`include "speed_neg_hs_test.sv" 
   	`include "token_in_test.sv" 
   	`include "debug_sof_test.sv" 
   	`include "token_out_ep1_test.sv" 
