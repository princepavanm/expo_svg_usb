interface sram_intf(input logic sram_clk, sram_rst);

  //Implement Modpot and clocking block here

endinterface:sram_intf
