//List of Include Files
  `include "usb_common.sv"
  `include "../reg/usb_reg_model.sv"
  `include "../reg/reg2wb_adapter.sv"

  `include "reset_intf.sv"
  `include "wb_intf.sv"
  `include "utmi_intf.sv"
  `include "sram_intf.sv"

  `include "reset_tx.sv"
  `include "reset_driver.sv"
  //`include "reset_sqr.sv"
  `include "reset_agent.sv"

  `include "wb_tx.sv"
  `include "wb_drv.sv"
  `include "wb_sqr.sv"
  `include "wb_cov.sv"
  `include "wb_mon.sv"
  `include "wb_agent.sv"

  `include "base_pkt.sv"

  `include "utmi_drv.sv"
  `include "utmi_sqr.sv"
  `include "utmi_cov.sv"
  `include "utmi_mon.sv"
  `include "utmi_agent.sv"

  `include "sram_tx.sv"
  `include "sram_drv.sv"
  `include "sram_sqr.sv"
  `include "sram_cov.sv"
  `include "sram_mon.sv"
  `include "sram_agent.sv"

  `include "virtual_sqr.sv"

// Sequence List
  `include "../seqs/wb_sequences/wb_seq_list.sv"
  `include "../seqs/utmi_sequences/utmi_seq_list.sv"
  `include "env.sv"
  `include "virtual_sequence.sv"

// Test List
  `include "../tests/test_list.sv"
