/* temp file for pushing purpose */
